CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
530 1210 3 110 10
176 79 1022 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 457 272
9437202 0
0
2 

2 

0
0
0
92
13 Logic Switch~
5 1309 149 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 20720 0
2 5V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5310 0 0
2
41384.6 0
0
13 Logic Switch~
5 1309 167 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 20720 0
2 5V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4318 0 0
2
41384.6 0
0
13 Logic Switch~
5 1309 186 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 20720 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3917 0 0
2
41384.6 0
0
13 Logic Switch~
5 1309 205 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 20720 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7930 0 0
2
41384.6 0
0
13 Logic Switch~
5 717 1538 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6128 0 0
2
41384.6 0
0
13 Logic Switch~
5 1082 265 0 1 11
0 15
0
0 0 21360 270
2 0V
-6 -21 8 -13
5 CLOCK
-18 -31 17 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7346 0 0
2
41384.6 0
0
13 Logic Switch~
5 33 950 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8577 0 0
2
5.89612e-315 0
0
13 Logic Switch~
5 1042 915 0 10 11
0 40 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3372 0 0
2
41384.6 1
0
13 Logic Switch~
5 1598 799 0 1 11
0 83
0
0 0 21360 90
2 0V
12 0 26 8
3 V12
9 -10 30 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3741 0 0
2
41384.6 2
0
13 Logic Switch~
5 1566 797 0 10 11
0 41 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V7
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5813 0 0
2
41384.6 3
0
13 Logic Switch~
5 577 792 0 10 11
0 44 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V6
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3213 0 0
2
41384.6 4
0
13 Logic Switch~
5 613 794 0 1 11
0 122
0
0 0 21360 90
2 0V
12 0 26 8
2 V1
12 -10 26 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3694 0 0
2
41384.6 5
0
5 4071~
219 84 951 0 3 22
0 16 16 18
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U18A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 17 0
1 U
4327 0 0
2
5.89612e-315 5.36716e-315
0
5 4049~
219 889 1598 0 2 22
0 20 19
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U17A
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 16 0
1 U
8800 0 0
2
5.89612e-315 5.37752e-315
0
5 4049~
219 968 1612 0 2 22
0 22 21
0
0 0 624 180
4 4049
-7 -24 21 -16
3 U9F
-5 -20 16 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 11 0
1 U
3406 0 0
2
5.89612e-315 5.38788e-315
0
5 4081~
219 925 1647 0 3 22
0 21 19 23
0
0 0 624 270
4 4081
-7 -24 21 -16
4 U16B
17 -4 45 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 15 0
1 U
6455 0 0
2
5.89612e-315 5.39306e-315
0
5 4081~
219 850 1648 0 3 22
0 21 20 24
0
0 0 624 270
4 4081
-7 -24 21 -16
4 U16A
17 -4 45 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 15 0
1 U
9319 0 0
2
5.89612e-315 5.39824e-315
0
14 Logic Display~
6 1012 1686 0 1 2
10 22
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 OF
-5 20 9 28
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3172 0 0
2
5.89612e-315 5.40342e-315
0
14 Logic Display~
6 923 1683 0 1 2
10 23
0
0 0 53872 180
6 100MEG
3 -16 45 -8
6 PERDEU
-19 20 23 28
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
38 0 0
2
5.89612e-315 5.4086e-315
0
14 Logic Display~
6 848 1682 0 1 2
31 24
0
0 0 53872 180
6 100MEG
3 -16 45 -8
6 GANHOU
-21 21 21 29
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
376 0 0
2
5.89612e-315 5.41378e-315
0
4 4585
219 848 1531 0 14 29
0 9 8 3 2 4 5 6 7 123
10 124 125 20 126
0
0 0 4848 270
4 4585
-14 -60 14 -52
7 COMPARA
-26 1 23 9
0
15 DVDD=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 2 7 10 14 1 9 11 4
6 5 12 3 13 15 2 7 10 14
1 9 11 4 6 5 12 3 13 0
65 0 0 512 1 0 0 0
1 U
6666 0 0
2
5.89612e-315 5.4371e-315
0
4 4008
219 865 1286 0 14 29
0 25 26 27 28 29 30 31 32 127
7 6 5 4 22
0
0 0 4848 270
4 4008
-14 -60 14 -52
7 SOMADOR
54 -7 103 1
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
9365 0 0
2
5.89612e-315 5.45264e-315
0
5 4027~
219 1097 1015 0 7 32
0 128 40 15 40 129 130 38
0
0 0 4720 0
4 4027
7 -60 35 -52
4 U13B
19 -61 47 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 13 0
1 U
3251 0 0
2
41384.6 6
0
5 4027~
219 1181 1015 0 7 32
0 131 40 38 40 132 133 37
0
0 0 4720 0
4 4027
7 -60 35 -52
4 U13A
19 -61 47 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 13 0
1 U
5481 0 0
2
41384.6 7
0
5 4027~
219 1349 1015 0 7 32
0 134 40 36 40 135 136 35
0
0 0 4720 0
4 4027
7 -60 35 -52
4 U12B
19 -61 47 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 12 0
1 U
7788 0 0
2
41384.6 8
0
5 4027~
219 1264 1015 0 7 32
0 137 40 37 40 138 139 36
0
0 0 4720 0
4 4027
7 -60 35 -52
4 U12A
19 -61 47 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 12 0
1 U
3273 0 0
2
41384.6 9
0
14 Logic Display~
6 1458 805 0 1 2
10 28
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3761 0 0
2
41384.6 10
0
14 Logic Display~
6 1433 805 0 1 2
10 27
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3226 0 0
2
41384.6 11
0
14 Logic Display~
6 1407 805 0 1 2
10 26
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4244 0 0
2
41384.6 12
0
14 Logic Display~
6 1381 805 0 1 2
10 25
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5225 0 0
2
41384.6 13
0
5 4049~
219 1128 900 0 2 22
0 38 28
0
0 0 624 90
4 4049
-7 -24 21 -16
3 U9D
16 -2 37 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 11 0
1 U
768 0 0
2
41384.6 14
0
5 4049~
219 1209 900 0 2 22
0 37 27
0
0 0 624 90
4 4049
-7 -24 21 -16
3 U9C
16 -2 37 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 11 0
1 U
5735 0 0
2
41384.6 15
0
5 4049~
219 1296 894 0 2 22
0 36 26
0
0 0 624 90
4 4049
-7 -24 21 -16
3 U9B
16 -2 37 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 11 0
1 U
5881 0 0
2
41384.6 16
0
5 4049~
219 1378 917 0 2 22
0 35 25
0
0 0 624 90
4 4049
-7 -24 21 -16
3 U9A
16 -2 37 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 11 0
1 U
3275 0 0
2
41384.6 17
0
5 7474~
219 218 1024 0 6 22
0 18 43 15 18 140 29
0
0 0 4720 0
4 7474
7 -60 35 -52
3 U8B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 10 0
1 U
4203 0 0
2
5.89612e-315 5.45523e-315
0
5 7474~
219 342 1024 0 6 22
0 18 29 15 18 141 30
0
0 0 4720 0
4 7474
7 -60 35 -52
3 U8A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 10 0
1 U
3440 0 0
2
5.89612e-315 5.45782e-315
0
5 7474~
219 472 1024 0 6 22
0 18 30 15 18 142 31
0
0 0 4720 0
4 7474
7 -60 35 -52
3 U7B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 9 0
1 U
9102 0 0
2
5.89612e-315 5.46041e-315
0
5 7474~
219 601 1024 0 6 22
0 18 31 15 42 143 32
0
0 0 4720 0
4 7474
7 -60 35 -52
3 U7A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 9 0
1 U
5586 0 0
2
5.89612e-315 5.463e-315
0
9 2-In XOR~
219 359 897 0 3 22
0 31 32 43
0
0 0 624 180
5 74F86
-18 -24 17 -16
3 U6A
-2 -25 19 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
525 0 0
2
5.89612e-315 5.46559e-315
0
14 Logic Display~
6 287 1242 0 1 2
10 29
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L1
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6206 0 0
2
5.89612e-315 5.46818e-315
0
14 Logic Display~
6 408 1243 0 1 2
10 30
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L2
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3418 0 0
2
5.89612e-315 5.47077e-315
0
14 Logic Display~
6 535 1243 0 1 2
10 31
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L3
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9312 0 0
2
5.89612e-315 5.47207e-315
0
14 Logic Display~
6 653 1243 0 1 2
10 32
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L4
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7419 0 0
2
5.89612e-315 5.47336e-315
0
2 +V
167 601 1048 0 1 3
0 42
0
0 0 53488 180
3 10V
8 -12 29 -4
3 V17
5 -22 26 -14
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
472 0 0
2
5.89612e-315 5.47466e-315
0
4 4514
219 1563 744 0 30 45
0 25 26 27 28 41 83 82 80 79
78 77 76 75 74 73 60 59 57 56
55 54 53 0 0 0 0 0 0 0
6
0
0 0 4848 90
4 4514
-14 -87 14 -79
2 U5
81 -6 95 2
0
16 DVDD=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 22 21 3 2 1 23 11 9 10
8 7 6 5 4 18 17 20 19 14
13 16 15 22 21 3 2 1 23 11
9 10 8 7 6 5 4 18 17 20
19 14 13 16 15 0
65 0 0 0 1 0 0 0
1 U
4714 0 0
2
41384.6 18
0
9 CC 7-Seg~
183 1182 174 0 18 19
10 52 51 50 49 48 47 46 45 144
2 2 2 2 2 2 2 2 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
7 COUNTER
-22 -57 27 -49
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
9386 0 0
2
41384.6 19
0
9 8-In NOR~
219 1120 488 0 9 19
0 82 79 78 76 75 74 73 60 72
0
0 0 624 90
4 4078
-7 -24 21 -16
2 A3
1 -2 15 6
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
7610 0 0
2
41384.6 20
0
9 8-In NOR~
219 1265 489 0 9 19
0 82 80 79 78 77 74 73 60 69
0
0 0 624 90
4 4078
-7 -24 21 -16
2 B3
0 -4 14 4
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
3482 0 0
2
41384.6 21
0
9 8-In NOR~
219 1411 489 0 9 19
0 82 80 78 77 76 75 74 73 70
0
0 0 624 90
4 4078
-7 -24 21 -16
2 C3
0 -2 14 6
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
3608 0 0
2
41384.6 22
0
9 8-In NOR~
219 1564 488 0 9 19
0 82 79 78 76 75 73 60 59 66
0
0 0 624 90
4 4078
-7 -24 21 -16
2 D1
1 -1 15 7
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
6397 0 0
2
41384.6 23
0
9 8-In NOR~
219 1685 486 0 9 19
0 82 79 75 73 59 56 145 146 81
0
0 0 624 90
4 4078
-7 -24 21 -16
2 E1
-1 -3 13 5
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 512 1 0 0 0
1 U
3967 0 0
2
41384.6 24
0
9 8-In NOR~
219 1758 487 0 9 19
0 82 77 76 75 73 60 59 54 64
0
0 0 624 90
4 4078
-7 -24 21 -16
2 F1
0 -2 14 6
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
8621 0 0
2
41384.6 25
0
9 8-In NOR~
219 1879 488 0 9 19
0 79 78 77 76 75 73 60 56 61
0
0 0 624 90
4 4078
-7 -24 21 -16
2 G3
1 -1 15 7
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
8901 0 0
2
41384.6 26
0
9 8-In NOR~
219 2001 488 0 9 19
0 59 57 56 55 54 53 147 148 62
0
0 0 624 90
4 4078
-7 -24 21 -16
4 dot1
-8 -1 20 7
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 512 1 0 0 0
1 U
7385 0 0
2
41384.6 27
0
9 Inverter~
13 1688 436 0 2 22
0 81 48
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11F
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
6519 0 0
2
41384.6 28
0
9 Inverter~
13 2003 439 0 2 22
0 62 45
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11E
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
552 0 0
2
41384.6 29
0
10 2-In NAND~
219 1160 426 0 3 22
0 72 71 52
0
0 0 624 90
4 7400
-7 -24 21 -16
3 U4D
19 -2 40 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
5551 0 0
2
41384.6 30
0
9 8-In NOR~
219 1193 488 0 9 19
0 59 56 55 53 149 150 151 152 71
0
0 0 624 90
4 4078
-7 -24 21 -16
2 A1
1 -1 15 7
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 512 1 0 0 0
1 U
8715 0 0
2
41384.6 31
0
10 2-In NAND~
219 1452 430 0 3 22
0 70 67 50
0
0 0 624 90
4 7400
-7 -24 21 -16
3 U4C
19 -2 40 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
9763 0 0
2
41384.6 32
0
9 8-In NOR~
219 1338 488 0 9 19
0 59 57 56 55 54 153 154 155 68
0
0 0 624 90
4 4078
-7 -24 21 -16
2 B1
-1 -2 13 6
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 512 1 0 0 0
1 U
8443 0 0
2
41384.6 33
0
10 2-In NAND~
219 1301 426 0 3 22
0 69 68 51
0
0 0 624 90
4 7400
-7 -24 21 -16
3 U4B
19 -2 40 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
3719 0 0
2
41384.6 34
0
9 8-In NOR~
219 1486 488 0 9 19
0 60 59 57 55 54 53 156 157 67
0
0 0 624 90
4 4078
-7 -24 21 -16
2 C1
-1 -2 13 6
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 512 1 0 0 0
1 U
8671 0 0
2
41384.6 35
0
9 4-In NOR~
219 1624 488 0 5 22
0 56 55 53 158 65
0
0 0 624 90
4 4002
-14 -24 14 -16
3 G1B
-5 0 16 8
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
11 typeDigital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 512 2 2 6 0
1 U
7168 0 0
2
41384.6 36
0
10 2-In NAND~
219 1597 428 0 3 22
0 66 65 49
0
0 0 624 90
4 7400
-7 -24 21 -16
3 U4A
19 -2 40 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
49 0 0
2
41384.6 37
0
9 Inverter~
13 1817 493 0 2 22
0 53 63
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11D
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
6536 0 0
2
41384.6 38
0
10 2-In NAND~
219 1789 428 0 3 22
0 64 63 47
0
0 0 624 90
4 7400
-7 -24 21 -16
3 U2D
19 -2 40 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3931 0 0
2
41384.6 39
0
10 2-In NAND~
219 1918 426 0 3 22
0 61 58 46
0
0 0 624 90
4 7400
-7 -24 21 -16
3 U2C
19 -2 40 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
4390 0 0
2
41384.6 40
0
9 4-In NOR~
219 1937 489 0 5 22
0 55 54 53 159 58
0
0 0 624 90
4 4002
-14 -24 14 -16
3 G1A
-3 -2 18 6
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
11 typeDigital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 512 2 1 6 0
1 U
3242 0 0
2
41384.6 41
0
9 4-In NOR~
219 948 494 0 5 22
0 94 93 92 160 97
0
0 0 624 90
4 4002
-14 -24 14 -16
2 G2
0 -2 14 6
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
11 typeDigital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 512 2 2 4 0
1 U
6760 0 0
2
41384.6 42
0
10 2-In NAND~
219 929 431 0 3 22
0 100 97 85
0
0 0 624 90
4 7400
-7 -24 21 -16
3 U2B
19 -2 40 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
5760 0 0
2
41384.6 43
0
10 2-In NAND~
219 800 433 0 3 22
0 103 102 86
0
0 0 624 90
4 7400
-7 -24 21 -16
3 U2A
19 -2 40 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3781 0 0
2
41384.6 44
0
9 Inverter~
13 828 498 0 2 22
0 92 102
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11C
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
8545 0 0
2
41384.6 45
0
10 2-In NAND~
219 608 433 0 3 22
0 105 104 88
0
0 0 624 90
4 7400
-7 -24 21 -16
3 U3D
19 -2 40 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
9739 0 0
2
41384.6 46
0
9 4-In NOR~
219 635 493 0 5 22
0 95 94 92 161 104
0
0 0 624 90
4 4002
-14 -24 14 -16
2 D2
-2 0 12 8
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
11 typeDigital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 512 2 1 4 0
1 U
388 0 0
2
41384.6 47
0
9 8-In NOR~
219 497 493 0 9 19
0 99 98 96 94 93 92 162 163 106
0
0 0 624 90
4 4078
-7 -24 21 -16
2 C2
-1 -2 13 6
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 512 1 0 0 0
1 U
4595 0 0
2
41384.6 48
0
10 2-In NAND~
219 312 431 0 3 22
0 108 107 90
0
0 0 624 90
4 7400
-7 -24 21 -16
3 U3C
19 -2 40 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3173 0 0
2
41384.6 49
0
9 8-In NOR~
219 349 493 0 9 19
0 98 96 95 94 93 164 165 166 107
0
0 0 624 90
4 4078
-7 -24 21 -16
2 B2
-1 -2 13 6
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 512 1 0 0 0
1 U
9261 0 0
2
41384.6 50
0
10 2-In NAND~
219 463 435 0 3 22
0 109 106 89
0
0 0 624 90
4 7400
-7 -24 21 -16
3 U3B
19 -2 40 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3494 0 0
2
41384.6 51
0
9 8-In NOR~
219 204 493 0 9 19
0 98 95 94 92 167 168 169 170 110
0
0 0 624 90
4 4078
-7 -24 21 -16
2 A2
1 -1 15 7
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 512 1 0 0 0
1 U
9101 0 0
2
41384.6 52
0
10 2-In NAND~
219 171 431 0 3 22
0 111 110 91
0
0 0 624 90
4 7400
-7 -24 21 -16
3 U3A
19 -2 40 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
358 0 0
2
41384.6 53
0
9 Inverter~
13 1014 444 0 2 22
0 101 84
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11B
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
3726 0 0
2
41384.6 54
0
9 Inverter~
13 699 441 0 2 22
0 120 87
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U10E
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
999 0 0
2
41384.6 55
0
9 8-In NOR~
219 1012 493 0 9 19
0 98 96 95 94 93 92 171 172 101
0
0 0 624 90
4 4078
-7 -24 21 -16
3 dot
-5 -1 16 7
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 512 1 0 0 0
1 U
8787 0 0
2
41384.6 56
0
9 8-In NOR~
219 890 493 0 9 19
0 118 117 116 115 114 112 99 95 100
0
0 0 624 90
4 4078
-7 -24 21 -16
1 G
4 -1 11 7
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
3348 0 0
2
41384.6 57
0
9 8-In NOR~
219 769 492 0 9 19
0 121 116 115 114 112 99 98 93 103
0
0 0 624 90
4 4078
-7 -24 21 -16
1 F
3 -2 10 6
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
3395 0 0
2
41384.6 58
0
9 8-In NOR~
219 696 491 0 9 19
0 121 118 114 112 98 95 173 174 120
0
0 0 624 90
4 4078
-7 -24 21 -16
1 E
2 -3 9 5
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 512 1 0 0 0
1 U
7740 0 0
2
41384.6 59
0
9 8-In NOR~
219 575 493 0 9 19
0 121 118 117 115 114 112 99 98 105
0
0 0 624 90
4 4078
-7 -24 21 -16
1 D
4 -1 11 7
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
6480 0 0
2
41384.6 60
0
9 8-In NOR~
219 422 494 0 9 19
0 121 119 117 116 115 114 113 112 109
0
0 0 624 90
4 4078
-7 -24 21 -16
1 C
3 -2 10 6
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
342 0 0
2
41384.6 61
0
9 8-In NOR~
219 276 494 0 9 19
0 121 119 118 117 116 113 112 99 108
0
0 0 624 90
4 4078
-7 -24 21 -16
1 B
3 -4 10 4
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
9953 0 0
2
41384.6 62
0
9 8-In NOR~
219 131 493 0 9 19
0 121 118 117 115 114 113 112 99 111
0
0 0 624 90
4 4078
-7 -24 21 -16
1 A
4 -2 11 6
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
361 0 0
2
41384.6 63
0
9 CC 7-Seg~
183 996 173 0 18 19
10 91 90 89 88 87 86 85 84 175
2 2 2 2 2 2 2 2 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
6 RANDOM
-17 -55 25 -47
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3343 0 0
2
41384.6 64
0
4 4514
219 574 749 0 30 45
0 29 30 31 32 44 122 121 119 118
117 116 115 114 113 112 99 98 96 95
94 93 92 0 0 0 0 0 0 0
9
0
0 0 4848 90
4 4514
-14 -87 14 -79
2 U1
81 -6 95 2
0
16 DVDD=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 22 21 3 2 1 23 11 9 10
8 7 6 5 4 18 17 20 19 14
13 16 15 22 21 3 2 1 23 11
9 10 8 7 6 5 4 18 17 20
19 14 13 16 15 0
65 0 0 0 1 0 0 0
1 U
7923 0 0
2
41384.6 65
0
299
1 4 2 0 0 12416 0 4 21 0 0 5
1321 205
2193 205
2193 1470
868 1470
868 1510
3 1 3 0 0 8320 0 21 3 0 0 5
877 1510
877 1456
2176 1456
2176 186
1321 186
5 13 4 0 0 4224 0 21 22 0 0 4
859 1510
859 1356
879 1356
879 1316
6 12 5 0 0 4224 0 21 22 0 0 4
850 1510
850 1347
870 1347
870 1316
7 11 6 0 0 4224 0 21 22 0 0 4
841 1510
841 1339
861 1339
861 1316
8 10 7 0 0 4224 0 21 22 0 0 4
832 1510
832 1331
852 1331
852 1316
2 1 8 0 0 12416 0 21 2 0 0 5
886 1510
886 1445
2162 1445
2162 167
1321 167
1 1 9 0 0 8320 0 1 21 0 0 5
1321 149
2148 149
2148 1435
895 1435
895 1510
1 10 10 0 0 4224 0 5 21 0 0 5
729 1538
782 1538
782 1502
805 1502
805 1510
0 0 11 0 0 0 0 0 0 0 0 2
921 1379
921 1379
0 0 12 0 0 0 0 0 0 0 0 2
884 1347
884 1347
0 0 13 0 0 0 0 0 0 0 0 2
879 1378
879 1378
0 0 14 0 0 0 0 0 0 0 0 2
870 1355
870 1355
0 1 15 0 0 8192 0 0 6 15 0 3
1007 826
1082 826
1082 277
3 0 15 0 0 12416 0 23 0 0 85 5
1073 988
1007 988
1007 826
140 826
140 1006
1 0 16 0 0 4096 0 7 0 0 17 2
45 950
60 950
1 2 16 0 0 8320 0 13 13 0 0 4
71 942
60 942
60 960
71 960
0 0 17 0 0 0 0 0 0 0 0 2
54 1032
54 1032
0 1 18 0 0 16512 0 0 38 38 0 8
157 951
157 1060
176 1060
176 1059
633 1059
633 956
601 956
601 961
2 2 19 0 0 8320 0 14 16 0 0 3
910 1598
914 1598
914 1625
0 1 20 0 0 4096 0 0 14 22 0 2
850 1598
874 1598
13 2 20 0 0 12416 0 21 17 0 0 4
850 1574
850 1598
839 1598
839 1626
1 0 21 0 0 4096 0 16 0 0 24 2
932 1625
932 1612
2 1 21 0 0 4224 0 15 17 0 0 3
953 1612
857 1612
857 1626
1 0 22 0 0 4096 0 15 0 0 26 2
989 1612
1012 1612
14 1 22 0 0 20608 0 22 18 0 0 8
897 1316
897 1368
949 1368
949 1373
1145 1373
1145 1578
1012 1578
1012 1672
3 1 23 0 0 4224 0 16 19 0 0 2
923 1670
923 1669
3 1 24 0 0 4224 0 17 20 0 0 2
848 1671
848 1668
0 1 25 0 0 8320 0 0 22 40 0 4
1513 828
1513 1185
897 1185
897 1252
0 2 26 0 0 8320 0 0 22 41 0 4
1522 835
1522 1174
888 1174
888 1252
0 3 27 0 0 8320 0 0 22 42 0 4
1531 839
1531 1164
879 1164
879 1252
0 4 28 0 0 8320 0 0 22 43 0 4
1540 844
1540 1154
870 1154
870 1252
5 0 29 0 0 8192 0 22 0 0 66 3
861 1252
861 1111
677 1111
6 0 30 0 0 8192 0 22 0 0 67 3
852 1252
852 1120
686 1120
7 0 31 0 0 8192 0 22 0 0 68 3
843 1252
843 1129
693 1129
8 0 32 0 0 8192 0 22 0 0 69 3
834 1252
834 1138
700 1138
0 0 33 0 0 0 0 0 0 0 0 2
59 999
59 999
3 1 18 0 0 0 0 13 37 0 0 3
117 951
472 951
472 961
0 0 34 0 0 4224 0 0 0 0 0 2
50 1045
50 1044
1 0 25 0 0 0 0 45 0 0 54 3
1513 775
1513 829
1381 829
2 0 26 0 0 0 0 45 0 0 46 3
1522 775
1522 835
1407 835
3 0 27 0 0 0 0 45 0 0 45 3
1531 775
1531 840
1433 840
4 0 28 0 0 0 0 45 0 0 44 3
1540 775
1540 845
1458 845
2 1 28 0 0 0 0 31 27 0 0 4
1131 882
1131 857
1458 857
1458 823
2 1 27 0 0 0 0 32 28 0 0 4
1212 882
1212 867
1433 867
1433 823
2 1 26 0 0 0 0 33 29 0 0 3
1299 876
1407 876
1407 823
1 7 35 0 0 4224 0 34 25 0 0 3
1381 935
1381 979
1373 979
1 0 36 0 0 4096 0 33 0 0 55 2
1299 912
1299 924
1 7 37 0 0 4224 0 32 24 0 0 3
1212 918
1212 979
1205 979
1 7 38 0 0 8320 0 31 23 0 0 4
1131 918
1130 918
1130 979
1121 979
3 0 36 0 0 4096 0 25 0 0 55 3
1325 988
1299 988
1299 978
3 0 37 0 0 0 0 26 0 0 49 3
1240 988
1212 988
1212 979
3 0 38 0 0 0 0 24 0 0 50 3
1157 988
1130 988
1130 977
1 2 25 0 0 0 0 30 34 0 0 2
1381 823
1381 899
0 7 36 0 0 4224 0 0 26 0 0 3
1299 918
1299 979
1288 979
0 0 39 0 0 0 0 0 0 0 0 2
1416 930
1416 930
2 0 40 0 0 4096 0 23 0 0 58 2
1073 979
1066 979
0 4 40 0 0 4096 0 0 23 64 0 3
1066 948
1066 997
1073 997
2 0 40 0 0 0 0 24 0 0 60 2
1157 979
1146 979
0 4 40 0 0 0 0 0 24 64 0 3
1146 948
1146 997
1157 997
2 0 40 0 0 0 0 26 0 0 62 2
1240 979
1232 979
0 4 40 0 0 0 0 0 26 64 0 3
1232 948
1232 997
1240 997
0 4 40 0 0 0 0 0 25 64 0 3
1317 979
1317 997
1325 997
1 2 40 0 0 8320 0 8 25 0 0 5
1042 927
1042 948
1317 948
1317 979
1325 979
5 1 41 0 0 4224 0 45 10 0 0 2
1567 775
1567 784
0 1 29 0 0 4224 0 0 92 73 0 5
287 1169
677 1169
677 860
524 860
524 780
0 2 30 0 0 8320 0 0 92 72 0 5
408 1178
686 1178
686 852
533 852
533 780
0 3 31 0 0 8320 0 0 92 71 0 5
535 1184
693 1184
693 846
542 846
542 780
0 4 32 0 0 8320 0 0 92 70 0 5
653 1192
700 1192
700 838
551 838
551 780
1 0 32 0 0 0 0 43 0 0 83 2
653 1229
653 988
1 0 31 0 0 0 0 42 0 0 86 2
535 1229
535 988
1 0 30 0 0 0 0 41 0 0 87 2
408 1229
408 988
1 0 29 0 0 0 0 40 0 0 88 2
287 1228
287 988
1 0 18 0 0 0 0 35 0 0 38 2
218 961
218 951
1 0 18 0 0 0 0 36 0 0 38 2
342 961
342 951
1 4 42 0 0 4224 0 44 38 0 0 2
601 1033
601 1036
4 0 18 0 0 0 0 35 0 0 19 2
218 1036
218 1059
4 0 18 0 0 0 0 36 0 0 19 2
342 1036
342 1059
4 0 18 0 0 0 0 37 0 0 19 2
472 1036
472 1059
3 0 15 0 0 0 0 37 0 0 85 3
448 1006
432 1006
432 1082
3 0 15 0 0 0 0 36 0 0 85 3
318 1006
306 1006
306 1082
3 2 43 0 0 4224 0 39 35 0 0 4
332 897
168 897
168 988
194 988
6 2 32 0 0 0 0 38 39 0 0 4
625 988
653 988
653 888
381 888
1 0 31 0 0 0 0 39 0 0 86 3
381 906
546 906
546 988
3 3 15 0 0 0 0 38 35 0 0 6
577 1006
567 1006
567 1082
140 1082
140 1006
194 1006
6 2 31 0 0 0 0 37 38 0 0 2
496 988
577 988
6 2 30 0 0 0 0 36 37 0 0 2
366 988
448 988
6 2 29 0 0 0 0 35 36 0 0 2
242 988
318 988
1 5 44 0 0 4224 0 11 92 0 0 2
578 779
578 780
2 8 45 0 0 8320 0 56 46 0 0 4
2006 421
2006 306
1203 306
1203 210
3 7 46 0 0 8320 0 67 46 0 0 4
1920 399
1920 301
1197 301
1197 210
3 6 47 0 0 8320 0 66 46 0 0 4
1791 401
1791 296
1191 296
1191 210
2 5 48 0 0 8320 0 55 46 0 0 4
1691 418
1691 291
1185 291
1185 210
3 4 49 0 0 8320 0 64 46 0 0 4
1599 401
1599 286
1179 286
1179 210
3 3 50 0 0 8320 0 59 46 0 0 4
1454 403
1454 388
1173 388
1173 210
3 2 51 0 0 12416 0 61 46 0 0 4
1303 399
1303 384
1167 384
1167 210
3 1 52 0 0 12416 0 57 46 0 0 4
1162 399
1162 384
1161 384
1161 210
22 3 53 0 0 8192 0 45 68 0 0 4
1495 711
1495 705
1948 705
1948 512
22 1 53 0 0 0 0 45 65 0 0 4
1495 711
1495 521
1820 521
1820 511
22 3 53 0 0 0 0 45 63 0 0 4
1495 711
1495 704
1635 704
1635 511
22 6 53 0 0 0 0 45 62 0 0 4
1495 711
1495 704
1506 704
1506 511
22 4 53 0 0 0 0 45 58 0 0 4
1495 711
1495 604
1195 604
1195 511
21 2 54 0 0 8192 0 45 68 0 0 4
1504 711
1504 705
1939 705
1939 512
21 8 54 0 0 0 0 45 52 0 0 4
1504 711
1504 703
1796 703
1796 510
21 5 54 0 0 0 0 45 62 0 0 4
1504 711
1504 704
1497 704
1497 511
21 5 54 0 0 0 0 45 60 0 0 4
1504 711
1504 614
1349 614
1349 511
20 1 55 0 0 8192 0 45 68 0 0 4
1513 711
1513 705
1930 705
1930 512
20 2 55 0 0 0 0 45 63 0 0 4
1513 711
1513 704
1626 704
1626 511
20 4 55 0 0 0 0 45 62 0 0 4
1513 711
1513 704
1488 704
1488 511
20 4 55 0 0 0 0 45 60 0 0 4
1513 711
1513 639
1340 639
1340 511
20 3 55 0 0 0 0 45 58 0 0 4
1513 711
1513 629
1186 629
1186 511
19 8 56 0 0 8192 0 45 53 0 0 4
1522 711
1522 704
1917 704
1917 511
19 6 56 0 0 0 0 45 51 0 0 4
1522 711
1522 707
1705 707
1705 509
19 1 56 0 0 0 0 45 63 0 0 4
1522 711
1522 704
1617 704
1617 511
19 3 56 0 0 0 0 45 60 0 0 4
1522 711
1522 634
1331 634
1331 511
19 2 56 0 0 0 0 45 58 0 0 4
1522 711
1522 619
1177 619
1177 511
22 6 53 0 0 8320 0 45 54 0 0 4
1495 711
1495 705
2021 705
2021 511
21 5 54 0 0 8320 0 45 54 0 0 4
1504 711
1504 705
2012 705
2012 511
20 4 55 0 0 8320 0 45 54 0 0 4
1513 711
1513 705
2003 705
2003 511
19 3 56 0 0 8320 0 45 54 0 0 4
1522 711
1522 705
1994 705
1994 511
18 2 57 0 0 8320 0 45 54 0 0 4
1531 711
1531 705
1985 705
1985 511
18 3 57 0 0 0 0 45 62 0 0 4
1531 711
1531 619
1479 619
1479 511
18 2 57 0 0 0 0 45 60 0 0 4
1531 711
1531 594
1322 594
1322 511
2 5 58 0 0 8320 0 67 68 0 0 4
1929 450
1929 455
1943 455
1943 456
17 1 59 0 0 8320 0 45 54 0 0 4
1540 711
1540 705
1976 705
1976 511
17 7 59 0 0 0 0 45 52 0 0 4
1540 711
1540 703
1787 703
1787 510
17 5 59 0 0 0 0 45 51 0 0 4
1540 711
1540 707
1696 707
1696 509
17 8 59 0 0 0 0 45 50 0 0 4
1540 711
1540 704
1602 704
1602 511
17 2 59 0 0 0 0 45 62 0 0 4
1540 711
1540 594
1470 594
1470 511
17 1 59 0 0 0 0 45 60 0 0 4
1540 711
1540 569
1313 569
1313 511
17 1 59 0 0 0 0 45 58 0 0 4
1540 711
1540 539
1168 539
1168 511
16 1 60 0 0 4096 0 45 62 0 0 4
1549 711
1549 539
1461 539
1461 511
9 1 61 0 0 8320 0 53 67 0 0 4
1885 455
1885 454
1911 454
1911 450
1 9 62 0 0 8320 0 56 54 0 0 3
2006 457
2007 457
2007 455
2 2 63 0 0 4224 0 65 66 0 0 3
1820 475
1820 452
1800 452
9 1 64 0 0 8320 0 52 66 0 0 3
1764 454
1764 452
1782 452
5 2 65 0 0 8320 0 63 64 0 0 3
1630 455
1630 452
1608 452
9 1 66 0 0 8320 0 50 64 0 0 3
1570 455
1570 452
1590 452
9 2 67 0 0 8320 0 62 59 0 0 3
1492 455
1492 454
1463 454
2 9 68 0 0 8320 0 61 60 0 0 3
1312 450
1312 455
1344 455
1 9 69 0 0 8320 0 61 48 0 0 3
1294 450
1294 456
1271 456
9 1 70 0 0 8320 0 49 59 0 0 3
1417 456
1417 454
1445 454
9 2 71 0 0 8320 0 58 57 0 0 3
1199 455
1199 450
1171 450
9 1 72 0 0 8320 0 47 57 0 0 4
1126 455
1126 456
1153 456
1153 450
16 7 60 0 0 8192 0 45 53 0 0 4
1549 711
1549 699
1908 699
1908 511
16 6 60 0 0 0 0 45 52 0 0 4
1549 711
1549 694
1778 694
1778 510
16 7 60 0 0 0 0 45 50 0 0 4
1549 711
1549 638
1593 638
1593 511
16 8 60 0 0 0 0 45 48 0 0 4
1549 711
1549 573
1303 573
1303 512
16 8 60 0 0 8320 0 45 47 0 0 4
1549 711
1549 544
1158 544
1158 511
15 6 73 0 0 8192 0 45 53 0 0 4
1558 711
1558 689
1899 689
1899 511
15 5 73 0 0 0 0 45 52 0 0 4
1558 711
1558 684
1769 684
1769 510
15 4 73 0 0 0 0 45 51 0 0 4
1558 711
1558 679
1687 679
1687 509
15 6 73 0 0 0 0 45 50 0 0 4
1558 711
1558 673
1584 673
1584 511
15 8 73 0 0 0 0 45 49 0 0 4
1558 711
1558 668
1449 668
1449 512
15 7 73 0 0 0 0 45 48 0 0 4
1558 711
1558 663
1294 663
1294 512
15 7 73 0 0 8320 0 45 47 0 0 4
1558 711
1558 659
1149 659
1149 511
14 7 74 0 0 12288 0 45 49 0 0 4
1567 711
1567 653
1440 653
1440 512
14 6 74 0 0 8192 0 45 48 0 0 4
1567 711
1567 648
1285 648
1285 512
14 6 74 0 0 8320 0 45 47 0 0 4
1567 711
1567 644
1140 644
1140 511
13 5 75 0 0 8192 0 45 53 0 0 4
1576 711
1576 649
1890 649
1890 511
13 4 75 0 0 0 0 45 52 0 0 4
1576 711
1576 644
1760 644
1760 510
13 3 75 0 0 0 0 45 51 0 0 4
1576 711
1576 639
1678 639
1678 509
13 5 75 0 0 0 0 45 50 0 0 4
1576 711
1576 633
1575 633
1575 511
13 6 75 0 0 0 0 45 49 0 0 4
1576 711
1576 628
1431 628
1431 512
13 5 75 0 0 8320 0 45 47 0 0 4
1576 711
1576 624
1131 624
1131 511
12 4 76 0 0 8192 0 45 53 0 0 4
1585 711
1585 629
1881 629
1881 511
12 3 76 0 0 0 0 45 52 0 0 4
1585 711
1585 624
1751 624
1751 510
12 4 76 0 0 0 0 45 50 0 0 4
1585 711
1585 618
1566 618
1566 511
12 5 76 0 0 0 0 45 49 0 0 4
1585 711
1585 613
1422 613
1422 512
12 4 76 0 0 8320 0 45 47 0 0 4
1585 711
1585 609
1122 609
1122 511
11 3 77 0 0 8192 0 45 53 0 0 4
1594 711
1594 614
1872 614
1872 511
11 2 77 0 0 0 0 45 52 0 0 4
1594 711
1594 609
1742 609
1742 510
11 4 77 0 0 0 0 45 49 0 0 4
1594 711
1594 603
1413 603
1413 512
11 5 77 0 0 8320 0 45 48 0 0 4
1594 711
1594 598
1276 598
1276 512
10 2 78 0 0 8192 0 45 53 0 0 4
1603 711
1603 599
1863 599
1863 511
10 3 78 0 0 0 0 45 50 0 0 4
1603 711
1603 593
1557 593
1557 511
10 3 78 0 0 0 0 45 49 0 0 4
1603 711
1603 588
1404 588
1404 512
10 4 78 0 0 8192 0 45 48 0 0 4
1603 711
1603 583
1267 583
1267 512
10 3 78 0 0 8320 0 45 47 0 0 4
1603 711
1603 579
1113 579
1113 511
9 1 79 0 0 8192 0 45 53 0 0 4
1612 711
1612 579
1854 579
1854 511
9 2 79 0 0 0 0 45 51 0 0 4
1612 711
1612 574
1669 574
1669 509
9 2 79 0 0 0 0 45 50 0 0 4
1612 711
1612 568
1548 568
1548 511
9 3 79 0 0 8192 0 45 48 0 0 4
1612 711
1612 563
1258 563
1258 512
9 2 79 0 0 8320 0 45 47 0 0 4
1612 711
1612 549
1104 549
1104 511
8 2 80 0 0 8192 0 45 49 0 0 4
1621 711
1621 558
1395 558
1395 512
8 2 80 0 0 8320 0 45 48 0 0 4
1621 711
1621 553
1249 553
1249 512
1 9 81 0 0 12416 0 55 51 0 0 4
1691 454
1691 455
1691 455
1691 453
7 1 82 0 0 4096 0 45 52 0 0 4
1630 711
1630 549
1733 549
1733 510
7 1 82 0 0 4096 0 45 51 0 0 4
1630 711
1630 544
1660 544
1660 509
7 1 82 0 0 4096 0 45 50 0 0 4
1630 711
1630 538
1539 538
1539 511
7 1 82 0 0 8192 0 45 49 0 0 4
1630 711
1630 533
1386 533
1386 512
7 1 82 0 0 8192 0 45 48 0 0 4
1630 711
1630 528
1240 528
1240 512
7 1 82 0 0 8320 0 45 47 0 0 4
1630 711
1630 524
1095 524
1095 511
6 1 83 0 0 8320 0 45 9 0 0 3
1585 781
1585 786
1599 786
2 8 84 0 0 4224 0 81 91 0 0 2
1017 426
1017 209
3 7 85 0 0 12416 0 70 91 0 0 4
931 404
931 389
1011 389
1011 209
3 6 86 0 0 8320 0 71 91 0 0 4
802 406
802 391
1005 391
1005 209
2 5 87 0 0 8320 0 82 91 0 0 4
702 423
702 408
999 408
999 209
3 4 88 0 0 8320 0 73 91 0 0 4
610 406
610 391
993 391
993 209
3 3 89 0 0 8320 0 78 91 0 0 4
465 408
465 301
987 301
987 209
3 2 90 0 0 8320 0 76 91 0 0 4
314 404
314 296
981 296
981 209
3 1 91 0 0 8320 0 80 91 0 0 4
173 404
173 291
975 291
975 209
22 3 92 0 0 8192 0 92 69 0 0 4
506 716
506 710
959 710
959 517
22 1 92 0 0 0 0 92 72 0 0 4
506 716
506 526
831 526
831 516
22 3 92 0 0 0 0 92 74 0 0 4
506 716
506 709
646 709
646 516
22 6 92 0 0 0 0 92 75 0 0 4
506 716
506 709
517 709
517 516
22 4 92 0 0 0 0 92 79 0 0 4
506 716
506 609
206 609
206 516
21 2 93 0 0 8192 0 92 69 0 0 4
515 716
515 710
950 710
950 517
21 8 93 0 0 0 0 92 85 0 0 4
515 716
515 708
807 708
807 515
21 5 93 0 0 0 0 92 75 0 0 4
515 716
515 709
508 709
508 516
21 5 93 0 0 0 0 92 77 0 0 4
515 716
515 619
360 619
360 516
20 1 94 0 0 8192 0 92 69 0 0 4
524 716
524 710
941 710
941 517
20 2 94 0 0 0 0 92 74 0 0 4
524 716
524 709
637 709
637 516
20 4 94 0 0 0 0 92 75 0 0 4
524 716
524 709
499 709
499 516
20 4 94 0 0 0 0 92 77 0 0 4
524 716
524 644
351 644
351 516
20 3 94 0 0 0 0 92 79 0 0 4
524 716
524 634
197 634
197 516
19 8 95 0 0 8192 0 92 84 0 0 4
533 716
533 709
928 709
928 516
19 6 95 0 0 0 0 92 86 0 0 4
533 716
533 712
716 712
716 514
19 1 95 0 0 0 0 92 74 0 0 4
533 716
533 709
628 709
628 516
19 3 95 0 0 0 0 92 77 0 0 4
533 716
533 639
342 639
342 516
19 2 95 0 0 0 0 92 79 0 0 4
533 716
533 624
188 624
188 516
22 6 92 0 0 8320 0 92 83 0 0 4
506 716
506 710
1032 710
1032 516
21 5 93 0 0 8320 0 92 83 0 0 4
515 716
515 710
1023 710
1023 516
20 4 94 0 0 8320 0 92 83 0 0 4
524 716
524 710
1014 710
1014 516
19 3 95 0 0 8320 0 92 83 0 0 4
533 716
533 710
1005 710
1005 516
18 2 96 0 0 8320 0 92 83 0 0 4
542 716
542 710
996 710
996 516
18 3 96 0 0 0 0 92 75 0 0 4
542 716
542 624
490 624
490 516
18 2 96 0 0 0 0 92 77 0 0 4
542 716
542 599
333 599
333 516
2 5 97 0 0 8320 0 70 69 0 0 4
940 455
940 460
954 460
954 461
17 1 98 0 0 8320 0 92 83 0 0 4
551 716
551 710
987 710
987 516
17 7 98 0 0 0 0 92 85 0 0 4
551 716
551 708
798 708
798 515
17 5 98 0 0 0 0 92 86 0 0 4
551 716
551 712
707 712
707 514
17 8 98 0 0 0 0 92 87 0 0 4
551 716
551 709
613 709
613 516
17 2 98 0 0 0 0 92 75 0 0 4
551 716
551 599
481 599
481 516
17 1 98 0 0 0 0 92 77 0 0 4
551 716
551 574
324 574
324 516
17 1 98 0 0 0 0 92 79 0 0 4
551 716
551 544
179 544
179 516
16 1 99 0 0 4096 0 92 75 0 0 4
560 716
560 544
472 544
472 516
9 1 100 0 0 8320 0 84 70 0 0 4
896 460
896 459
922 459
922 455
1 9 101 0 0 8320 0 81 83 0 0 3
1017 462
1018 462
1018 460
2 2 102 0 0 4224 0 72 71 0 0 3
831 480
831 457
811 457
9 1 103 0 0 8320 0 85 71 0 0 3
775 459
775 457
793 457
5 2 104 0 0 8320 0 74 73 0 0 3
641 460
641 457
619 457
9 1 105 0 0 8320 0 87 73 0 0 3
581 460
581 457
601 457
9 2 106 0 0 8320 0 75 78 0 0 3
503 460
503 459
474 459
2 9 107 0 0 8320 0 76 77 0 0 3
323 455
323 460
355 460
1 9 108 0 0 8320 0 76 89 0 0 3
305 455
305 461
282 461
9 1 109 0 0 8320 0 88 78 0 0 3
428 461
428 459
456 459
9 2 110 0 0 8320 0 79 80 0 0 3
210 460
210 455
182 455
9 1 111 0 0 8320 0 90 80 0 0 4
137 460
137 461
164 461
164 455
16 7 99 0 0 8192 0 92 84 0 0 4
560 716
560 704
919 704
919 516
16 6 99 0 0 0 0 92 85 0 0 4
560 716
560 699
789 699
789 515
16 7 99 0 0 0 0 92 87 0 0 4
560 716
560 643
604 643
604 516
16 8 99 0 0 0 0 92 89 0 0 4
560 716
560 578
314 578
314 517
16 8 99 0 0 8320 0 92 90 0 0 4
560 716
560 549
169 549
169 516
15 6 112 0 0 8192 0 92 84 0 0 4
569 716
569 694
910 694
910 516
15 5 112 0 0 0 0 92 85 0 0 4
569 716
569 689
780 689
780 515
15 4 112 0 0 0 0 92 86 0 0 4
569 716
569 684
698 684
698 514
15 6 112 0 0 0 0 92 87 0 0 4
569 716
569 678
595 678
595 516
15 8 112 0 0 0 0 92 88 0 0 4
569 716
569 673
460 673
460 517
15 7 112 0 0 0 0 92 89 0 0 4
569 716
569 668
305 668
305 517
15 7 112 0 0 8320 0 92 90 0 0 4
569 716
569 664
160 664
160 516
14 7 113 0 0 12288 0 92 88 0 0 4
578 716
578 658
451 658
451 517
14 6 113 0 0 8192 0 92 89 0 0 4
578 716
578 653
296 653
296 517
14 6 113 0 0 8320 0 92 90 0 0 4
578 716
578 649
151 649
151 516
13 5 114 0 0 8192 0 92 84 0 0 4
587 716
587 654
901 654
901 516
13 4 114 0 0 0 0 92 85 0 0 4
587 716
587 649
771 649
771 515
13 3 114 0 0 0 0 92 86 0 0 4
587 716
587 644
689 644
689 514
13 5 114 0 0 0 0 92 87 0 0 4
587 716
587 638
586 638
586 516
13 6 114 0 0 0 0 92 88 0 0 4
587 716
587 633
442 633
442 517
13 5 114 0 0 8320 0 92 90 0 0 4
587 716
587 629
142 629
142 516
12 4 115 0 0 8192 0 92 84 0 0 4
596 716
596 634
892 634
892 516
12 3 115 0 0 0 0 92 85 0 0 4
596 716
596 629
762 629
762 515
12 4 115 0 0 0 0 92 87 0 0 4
596 716
596 623
577 623
577 516
12 5 115 0 0 0 0 92 88 0 0 4
596 716
596 618
433 618
433 517
12 4 115 0 0 8320 0 92 90 0 0 4
596 716
596 614
133 614
133 516
11 3 116 0 0 8192 0 92 84 0 0 4
605 716
605 619
883 619
883 516
11 2 116 0 0 0 0 92 85 0 0 4
605 716
605 614
753 614
753 515
11 4 116 0 0 0 0 92 88 0 0 4
605 716
605 608
424 608
424 517
11 5 116 0 0 8320 0 92 89 0 0 4
605 716
605 603
287 603
287 517
10 2 117 0 0 8192 0 92 84 0 0 4
614 716
614 604
874 604
874 516
10 3 117 0 0 0 0 92 87 0 0 4
614 716
614 598
568 598
568 516
10 3 117 0 0 0 0 92 88 0 0 4
614 716
614 593
415 593
415 517
10 4 117 0 0 8192 0 92 89 0 0 4
614 716
614 588
278 588
278 517
10 3 117 0 0 8320 0 92 90 0 0 4
614 716
614 584
124 584
124 516
9 1 118 0 0 8192 0 92 84 0 0 4
623 716
623 584
865 584
865 516
9 2 118 0 0 0 0 92 86 0 0 4
623 716
623 579
680 579
680 514
9 2 118 0 0 0 0 92 87 0 0 4
623 716
623 573
559 573
559 516
9 3 118 0 0 8192 0 92 89 0 0 4
623 716
623 568
269 568
269 517
9 2 118 0 0 8320 0 92 90 0 0 4
623 716
623 554
115 554
115 516
8 2 119 0 0 8192 0 92 88 0 0 4
632 716
632 563
406 563
406 517
8 2 119 0 0 8320 0 92 89 0 0 4
632 716
632 558
260 558
260 517
1 9 120 0 0 12416 0 82 86 0 0 4
702 459
702 460
702 460
702 458
7 1 121 0 0 4096 0 92 85 0 0 4
641 716
641 554
744 554
744 515
7 1 121 0 0 4096 0 92 86 0 0 4
641 716
641 549
671 549
671 514
7 1 121 0 0 4096 0 92 87 0 0 4
641 716
641 543
550 543
550 516
7 1 121 0 0 8192 0 92 88 0 0 4
641 716
641 538
397 538
397 517
7 1 121 0 0 8192 0 92 89 0 0 4
641 716
641 533
251 533
251 517
7 1 121 0 0 8320 0 92 90 0 0 4
641 716
641 529
106 529
106 516
6 1 122 0 0 4224 0 92 12 0 0 4
596 786
605 786
605 781
614 781
6
-32 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
1232 147 1266 201
1239 154 1258 190
1 =
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1277 134 1298 155
1283 141 1291 156
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1276 171 1299 192
1283 178 1291 193
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1275 191 1300 212
1283 198 1291 213
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1274 153 1301 174
1283 159 1291 174
1 4
-32 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
1067 145 1112 203
1079 155 1099 193
1 +
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
